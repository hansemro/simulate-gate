
* set gnd and power
.PARAM vdd = 1.8
Vgnd VGND 0 0
Vdd VPWR VGND vdd

* create a pulse for A 
Va A VGND pulse(0 1.8 1n 10p 10p 1n 2n)

Vb B VGND pulse(0 1.8 1.5n 10p 10p 1n 2n)

* setup the transient analysis
.tran 10p 3n 0

* fall delay
.meas TRAN fall_delay
    + TRIG V(A) VAL='0.5*vdd' TD=0 FALL=1
    + TARG V(Y) VAL='0.5*vdd' TD=0 RISE=1

* rise delay
.meas TRAN rise_delay
    + TRIG V(B) VAL='0.5*vdd' TD=0 RISE=1
    + TARG V(Y) VAL='0.5*vdd' TD=0 FALL=1

* rise time
.meas TRAN rise_time
    + TRIG V(Y) VAL='0.2*vdd' TD=0 RISE=1
    + TARG V(Y) VAL='0.8*vdd' TD=0 RISE=1

* fall time
.meas TRAN fall_time
    + TRIG V(Y) VAL='0.8*vdd' TD=0 FALL=1
    + TARG V(Y) VAL='0.2*vdd' TD=0 FALL=1

.control
run
set color0 = white
set color1 = black
plot A B Y
.endc

.end
